`timescale 1ns/1ps

module display_480p_tb();
	logic clk, rst, hsync, vsync, de, frame, line;
	logic [15:0] screen_x, screen_y;
//	display_480p ()
//	initial begin
//		display_item item;
//		repeat (width) begin
//			@(posedge clk) line_signal: assert (line);
//		end
//	end
endmodule


//class display_item;
//	logic clk, rst, hsync, vsync, de, frame, line;
//	logic [15:0] screen_x, screen_y;
//	
//endclass
